Fuzz Tone

.include fuzztone.mod

* calculate bias at minimum attack
.param att=0.01
.param vol=0.99

* original values from patent
.param r19=10k
.param r26=1.5k
.param r35=10k

X1 in out fuzztone att=att vol=vol r19=r19 r26=r26 r35=r35

.param amp=1

Vin in 0 sin(0 {amp} 440 0 0)

.control

let targ_v2 = -1.5
let best_v2 = 100
let best_v2err = 100

let targ_v7 = -3
let best_v7 = 100
let best_v7err = 100

let targ_v9 = -2.5
let best_v9 = 100
let best_v9err = 100


let start_r19 = 100
let stop_r19 = 20k
let delta_r19 = 100
let r19_act = start_r19
let best_r19 = 10k

let start_r26 = 100
let stop_r26 = 10k
let delta_r26 = 100
let r26_act = start_r26
let best_r26 = 1.5k

let start_r35 = 100
let stop_r35 = 20k
let delta_r35 = 100
let r35_act = start_r35
let best_r35 = 10k


* loop
while r19_act < stop_r19

alterparam r19 = $&r19_act
reset
op

let v2err = abs(v(x1.2)-targ_v2)
if v2err le best_v2err
let best_v2 = v(x1.2)
let best_v2err = v2err
let best_r19 = r19_act
end

let r19_act = r19_act + delta_r19
end


* loop
while r26_act < stop_r26

alterparam r19 = $&best_r19
alterparam r26 = $&r26_act
reset
op

let v7err = abs(v(x1.7)-targ_v7)
if v7err le best_v7err
let best_v7 = v(x1.7)
let best_v7err = v7err
let best_r26 = r26_act
end

let r26_act = r26_act + delta_r26
end


* loop
while r35_act < stop_r35

alterparam r19 = $&best_r19
alterparam r26 = $&best_r26
alterparam r35 = $&r35_act
reset
op

let v9err = abs(v(x1.9)-targ_v9)
if v9err le best_v9err
let best_v9 = v(x1.9)
let best_v9err = v9err
let best_r35 = r35_act
end

let r35_act = r35_act + delta_r35
end


print best_r19
print best_r26
print best_r35


alterparam r19 = $&best_r19
alterparam r26 = $&best_r26
alterparam r35 = $&best_r35
reset
op

let best_v2 = v(x1.2)
let best_v7 = v(x1.7)
let best_v9 = v(x1.9)

tran 22.675u 0.009

print targ_v2 best_v2
print targ_v7 best_v7
print targ_v9 best_v9

.endc

.end
